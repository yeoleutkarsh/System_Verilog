
interface intf;
  
  logic a;
  logic b;
  logic sum;
  logic carry;
  
  // It also contain clocking block
  // and modport -> to bundle the signal.
endinterface
