
interface intf ( input logic clk, rst );
    logic [3:0] in1;
    logic [3:0] in2;
    logic [4:0] out; 
endinterface
